module Instruction_Memory(
    input CLK,
    input RST,
    input [31:0]address,
    output reg [31:0] instruction,
);



endmodule