
module HazardDetector(
    input HD_instruction,
    input [1:0] HD_IDEX_memread,
    input [2:0]HD_Rx_a_IDEX,
    input [2:0]HD_Ry_a_IDEX,
    output PCWrite,
    output IFIDWrite,
    output addBubble
    
    );
    
    if( HD_IDEX_memread[1:0] == )
    
    
    
endmodule
